`timescale 1ns/1ps
module top_test;
  reg clk;
  reg rst;
  reg PB0;
  reg PB1;
  reg PB2;
  reg[7:0]SW;
  wire [3:0]AN;
  wire [7:0]LED;
  wire [6:0]seg;
  TOP_ALU top_alu(clk,rst,PB0,PB1,PB2,SW,LED,AN,seg);
  integer i;
  initial begin
  clk=0; rst=1; PB0=0; PB1=0; PB2=0; SW=0;
  #1 rst = 0;
  #5000000 PB0 = 1 ; SW = 255;
  #10000000 PB0 = 0;
  #5000000 PB1=1; SW=15;
  #10000000 PB1=0;
  SW=0;
  for(i=0;i<7;i=i+1)
  begin
    #5000000 PB2=1; SW=SW+1;
    #10000000 PB2=0;
  end
end
always #10 clk= ~clk;
endmodule
  initial begin
  clk = 0;
  forever #10 clk = ~clk;
  end
  initial begin
  $monitor($time,,,,"rst=%b , PB0=%b , PB1=%b , PB2=%b , SW=%b , LED=%b , seg=%b  ",rst,PB0,PB1,PB2,SW,LED,AN,seg);
  SW=8'b00110010;
  #1000000;
  PB0 =1;
  #2000;
  PB0 = 0;
  #1000;
  PB0 =1;
  #3000; 
  PB0 = 0;
  #1000;
  PB0 =1;
  #4000;
  PB0 = 0;
  #1000;
  PB0 =1;
  #3000; 
  PB0 = 0;
  #1000;
  PB0 =1; 
  #10000000; 
  PB0 = 0;
  #1000;
  PB0 =1;
  #2000;
  PB0 = 0;
  #1000;
  PB0 =1;
  #3000; 
  PB0 = 0;
  #5000000;
  SW=8'b01001011;
  #5000000;
  PB1 = 0;
  #1000;
  PB1 =1;
  #2000;
  PB1 = 0;
  #1000;
  PB1 =1;
  #3000; 
  PB1 = 0;
  #1000;
  PB1 =1;
  #4000;
  PB1 = 0;
  #1000;
  PB1 =1;
  #3000; 
  PB1 = 0;
  #1000;
  PB1 =1; 
  #10000000; 
  PB1 = 0;
  #1000;
  PB1 =1;
  #2000;
  PB1 = 0;
  #1000;
  PB1 =1;
  #3000; 
  PB1 = 0;
  #5000000;
  SW=8'b00000001;
  #5000000;
  PB2 = 0;
  #1000;
  PB2 =1;
  #2000;
  PB2 = 0;
  #1000;
  PB2 =1;
  #3000; 
  PB2 = 0;
  #1000;
  PB2 =1;
  #4000;
  PB2 = 0;
  #1000;
  PB2 =1;
  #3000; 
  PB2 = 0;
  #1000;
  PB2 =1; 
  #10000000; 
  PB2 = 0;
  #1000;
  PB2 =1;
  #2000;
  PB2 = 0;
  #1000;
  PB2 =1;
  #3000; 
  PB2 = 0;
  end
